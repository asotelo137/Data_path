/****************************************************************************
 * if_df_buffer.sv
 ****************************************************************************/

/**
 * Module: if_df_buffer
 * 
 * TODO: Add module documentation
 */
module if_df_buffer;


endmodule


